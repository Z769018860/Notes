`timescale 10 ns / 1 ns

`define DATA_WIDTH 32
`define AND 3'b000
`define OR 3'b001
`define ADD 3'b010
`define SUB 3'b110
`define SLT 3'b111
`define todo 1
`define UNDEFINED 0

module alu(
	input [`DATA_WIDTH - 1:0] A,
	input [`DATA_WIDTH - 1:0] B,
	input [2:0] ALUop,
	output Overflow,
	output CarryOut,
	output Zero,
	output [`DATA_WIDTH - 1:0] Result
);

    wire [`DATA_WIDTH-1:0] Chooser;
    assign Chooesr=
//Zero
	assign Zero=({Result}==0);

    assign {CarryOut,Reuslt}=
        &&
endmodule
